
/* ****************************************************************************
  This Source Code Form is subject to the terms of the
  Open Hardware Description License, v. 1.0. If a copy
  of the OHDL was not distributed with this file, You
  can obtain one at http://juliusbaxter.net/ohdl/ohdl.txt
  
  Copyright (C) 2019 Stefan Huemer <stefan@huemer.tech>
  
***************************************************************************** */

`define ASCII_WIDTH ( 7 )

`define ASCII_LF    ( 10 )
`define ASCII_SPACE ( 32 )

`define ASCII_0     ( 48 )
