
/* ****************************************************************************
  This Source Code Form is subject to the terms of the
  Open Hardware Description License, v. 1.0. If a copy
  of the OHDL was not distributed with this file, You
  can obtain one at http://juliusbaxter.net/ohdl/ohdl.txt
  
  Copyright (C) 2019 Stefan Huemer <stefan@huemer.tech>
  
***************************************************************************** */

//~ parameter MEM_SIZE = 4194304 + 1;
//~ parameter MEM_SIZE = 14194304 + 1;
//~ parameter MEM_SIZE = ( 17 * 262144 ) + 1;

//~ `define MEM_SIZE ( ( 17 * 262144 ) + 1 )

//`define MEM_SIZE ( (3 * 25048) + 1 )
//`define MEM_SIZE ( (3 * 2048) + 1 )

`define MEM_SIZE ( 100192 )

