
/* ****************************************************************************
  This Source Code Form is subject to the terms of the
  Open Hardware Description License, v. 1.0. If a copy
  of the OHDL was not distributed with this file, You
  can obtain one at http://juliusbaxter.net/ohdl/ohdl.txt
  
  Copyright (C) 2019 Stefan Huemer <stefan@huemer.tech>
  
***************************************************************************** */

`define N0_ARCH ( `RV32I )
`define N1_ARCH ( `RV32IM )
`define N2_ARCH  ( 1'b1 )
`define N3_ARCH  ( 1'b1 )
`define N4_ARCH  ( 1'b1 )
`define N5_ARCH  ( 1'b1 )
`define N6_ARCH  ( 1'b1 )
`define N7_ARCH  ( 1'b1 )
`define N8_ARCH  ( 1'b1 )
`define N9_ARCH  ( 1'b1 )
`define N10_ARCH ( 1'b1 )
`define N11_ARCH ( 1'b1 )
`define N12_ARCH ( 1'b1 )
`define N13_ARCH ( 1'b1 )
`define N14_ARCH ( 1'b1 )
`define N15_ARCH ( 1'b1 )
`define N16_ARCH ( 1'b1 )
`define N17_ARCH ( 1'b1 )
`define N18_ARCH ( 1'b1 )
`define N19_ARCH ( 1'b1 )
`define N20_ARCH ( 1'b1 )
`define N21_ARCH ( 1'b1 )
`define N22_ARCH ( 1'b1 )
`define N23_ARCH ( 1'b1 )
`define N24_ARCH ( 1'b1 )
`define N25_ARCH ( 1'b1 )
`define N26_ARCH ( 1'b1 )
`define N27_ARCH ( 1'b1 )
`define N28_ARCH ( 1'b1 )
`define N29_ARCH ( 1'b1 )
