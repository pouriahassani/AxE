
/* ****************************************************************************
  This Source Code Form is subject to the terms of the
  Open Hardware Description License, v. 1.0. If a copy
  of the OHDL was not distributed with this file, You
  can obtain one at http://juliusbaxter.net/ohdl/ohdl.txt
  
  Copyright (C) 2019 Stefan Huemer <stefan@huemer.tech>
  
***************************************************************************** */
// sobel 8x8 needs this much memory!!!
`define MEM_SIZE ( 268435455 )
// `define MEM_SIZE ( 2048 )
// `define MEM_SIZE ( 36880 )

`define MEM_PATH ( "/home/user/soc_frame/mem.hex" )
