`define PATH_IF_AXI_LIGHT ( "../../../rtl/interfaces/if_axi_light.sv" )

`define PATH_AXI_DETECTOR ( "../../../rtl/axi_detector/axi_detector.sv" )

`define PATH_PICORV32 ( "../../../rtl/pico/picorv32.v" )

`define PATH_PICORV32_IF_WRAPPER_CADENCE ( "../../../rtl/pico/picorv32_if_wrapper_cadence.sv" )

`define PATH_MEMORY_ASIC_MEMORY_LATCH1 ( "../../../rtl/memory_asic/memory_latch1.sv" )
`define PATH_MEMORY_ASIC_LATCH_REGISTER_FILE ( "../../../rtl/memory_asic/latch_register_file.sv" )
`define PATH_MEMORY_ASIC_LATCH_REGISTER_FILE_WRAPPER ( "../../../rtl/memory_asic/latch_register_file_wrapper.sv" )
`define PATH_MEMORY_ASIC_CLUSTER_CLOCK_GATING ( "../../../rtl/memory_asic/cluster_clock_gating.sv" )

`define PATH_PICORV32_IF_WRAPPER ( "../../../rtl/pico/picorv32_if_wrapper.sv" )

`define PATH_MEMORY_MEM_PACKER ( "../../../rtl/memory/memory_mem_packer.sv" )

`define PATH_DEBUGGER ( "../../../rtl/debugger/debugger.sv" )
